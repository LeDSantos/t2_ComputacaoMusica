BZh91AY&SYG,T# [D߀Ryg����������`=�}B+�   ;s�x���g\  �	�ۛ]iM��@)����\5[1KZ�leJIT�:�+q]��a��2(Ln	�l2����N�)"�Gc �<� !�
(T����� �  � dS�%T��i�0  �M08ɓF!���`��i�5?F�$Pdb4  ��A�F� ���Tߪ���?'�LMM�ަ�� @�4L�ț*zOS�~�DzM=O(h4�Mn��󢈧�(ZJ
b�E �  T�2(����?�y�D��(P�5�5�����#b���CSYMx\�ND�}6����c�:4~������_u����X|�')�eo!EΘ�M���̨�cX*I(�qZePlR�H$�9{Gh��q/s� ���Y��4�r��ǎ6�{�N1MB?�0V���������z�Pa�/Yݛ0t��q���!N�U�hÅ4
��}�D\>1TJDP$�:b"��h�PU�N�O_ۊ[9���k[��g)�l8V�I����ǧ�]��u�����x�����1�
0��*^]۷�����R$�u��z�c�mM�U��Mc)��z�B���V䵕*ZF�k'�Ա�#�����ldIumRT�8�+�`��8�D|^�6O�¾%W�4��ȑ�V@������U�S���ɺ��{*�V)ié�Ui�qeѿB�Q^��Ѣ�ّ��髣6��
�:*�c�d�v׀�좽u�ۢ�۽�sw���ö�g���8ۢf�/h�aՖL���P���d�,�+��x���U��6����1vê1�3Y�nÔ�j��<�t��X7R����M�R��!�E1W����(e�B��1��X��l[TE�fZ�b�6��HB�AQm#/4e��m*�pe�	�.[��p���˻Ӈ)ʥb�㻎����Y����T�R,�e+aٛ�F�8oP�&V�#1n��[�&����jn�E�X��sAC&f��{`ݷD��k.�lz�WHe�;���ٰ���j�R#kV��]*�~vA����O�����jeJ�s�������WB0�̬�B��E�3�'P�)b��*�\��ݵ�҇��dkf��8M{/����&qۿ=9���=��Ex�cM�i���*�h�1R11�afS��n��*��X����[n��Z�U���x�O3e�=�A.��GPh�ot��j�h�w��k�V�f]߼����*cp��V�4���ep��i��
���gBF�!�Ɲ\s�^�t,p^�Y"���7�X;���.�m������6��Z>X���?�F?�?�~W��6Lf:�a'�۳�.��I�ꬾ�7���0!a�-�,4�o�=�;;z�V��E�S��٭;8c@��(��hu�a�N�363^<����������?W�i��\�\�[
,-X�Kvՙs��sn����i�ic��f�f�Y�]���P���U*�9�i�Vڿn��u�R�[e���tn`�E����P�˴����b����W.~�g��?O��#O���HW}�"w��-�^F�so�t���GV�=�"׵Wtw��	eA��r�
N:��T[k{���|c(\�Q�{���5Y�����\��M����0,g��i�M@a��e��'+2�K�l�e��Q���4�\욑�Ʋ�M-W1T�em4s2ڱ����!��b��)M�1��щ��ōI_~�Gq{�E5��3cbQGW��#-�[,�u]6�r�lB7%��DR��/�}k��ٳ��bwv��-�H�C"I��r�6@�
B�]6!n��%��B��j?Q�w[���6�,�0��m�������Raf�gQ�F5��Wf��h�˫6���.�\K+˖���ڥX˸�ˉM�J���%���̦�kL:�Mk0��И��F��s8�X4�pC]Y��fYb��{�~>�Mu�ֺK^ҵ�4D��q���r�RJ�;}Z�P�ky�|zqzk7�4zS���ņ��~ϝ��9 �7������������L�D�����E����c613?��hҤ�dS��B��Y	�V�ʆ�Y�-۽�HYTFV�i�s��ݾ]Zl�N2�>G��J�����LR�Z�!g�6�UX(��ԑ�XD˨RJ�Z�ei�p48�K�e6I��R�H�j��i�)]a��ǈ�最�X-�Ӽ���R�7�Q*��Q�["�[��{��cqa��P�>wSՑ��U�v��^;/��^"af�hw�ر�TNF倆K�h-���cl6��K�E*[qKtY��էmإ)F��;k0q�=F]:b%��'���%mꮻ�Gg^�;d������[u:5OSz񌻻����6$b�d�U�}��tO�4��1#;�f�c�n��dV�i9v��c��P)������F�4v�u%��PDu{,��p߳�tY�ͳ�>a��fN-5x�Xl(�Y�5�� x�/A	[�x�l\vF�W7�U�\����y�iŷ���%��oL�fc�o3I*�����QZ��T闘ڙe9�ٷ)��P+�ũ�+k��L�}$ճf����O�D������D�c��/����F�v�ަ�p�St##7�)�����]�n���T� ^)��c[�:ڮq.պ۵�V����ۓl��������׋Q��պ7Qt�m��ȳw�{�=��Ⱦbh$�gz�b��:1��Vm[��a��l�m����Q`9�4^�(sq��Eڨ$D�Y*/�hoFZb��Tah�%%�A^�V��[N�A�D�N�:)�ь�3^�s���츟�_�$=y����g�z*�\IW��uǋnǝ��q¼ɽ�H�^�  v۟E�f���9���E��j��^h����@��� �D]�x9K84�{oz�TE��V:	�Lx�2�;�芢Y�2%^taⵥ7���{���1T߷�оXC����B,4hJh��lG&@�#Gg��Ht��	�Aug'ɠn��N���jc��V+c�^�&8_��4��m}� M����ɘX�����j����+�U����Ӫ�ŝg��Ы�Z���w���p�K��o3eȫs�{�bæge�qСݺ�u�l�Z�fůӰ���&/-�?%�'V���0A�g�g(�(e�_���hُ͎%^�mF��@2���"���ǻp3�z�Mz;�۶�SYp�7-w/�b�J�{�LU܋��v����� u���>�{aQp�r-M9��v��r<{���~ �D?���>:(�I$R  ��!��9ڗ�ؖm%����a-��
��X�	Ub�B���T�����h ���� �ȅY�e�s *�1\_s.q��b5��l��f_��~n$Z� �����@ ��Ә���{�'��`�Dx_���LȒY�Or�\eڳ[o���N�O<(������q��
j����<H��F��u)����:(���@�Z�J��\z�]�
t �s�C�gRl��Y`�DM �/�mC�@ހ�A�?�g�/WDxy�H]�Dh�+#�"|�\4��3�^��Ȑ>H�L���j?! F�`��B��$5�9�J�)�|�O�Q���^��j��ڡO���&	�:v�vb�j�������'��<ᢁQ�"$N��gm�0�G�Z/�C|��<�xxF#V|Û{][nɁ9�,��3��m��t��5�Ub[c��9����,L<G������:C���0O��b�n?g�c��F��2c9ظfgii��ny�V��z!����v���H �V5tt*ݡC�k��P��a�V����ʜ�	 ��U2B��HMYh�k�b�s\n�	Q�����C_� ;���!�Z���,�C����h@D�=R��^�]�{�ru�+�/
�Ǳ��d��G�\�D0����޾���C=Hxh>�B  ,qc�2Mg}RI=���R�ru�Պ��v������ϥ��6��nV�e��Pv�o��i[�*�n��۝�:�]����Q�5KW��F�.�����͹5�+hl���c�/��H A҈
B��=A��^^�˜�Y��&9�?�? /������u�����#﯃>M�S; �}�%�D�W���s��+ �.=.s_��w��ʈ� ��!��X���Ś�[���y��=�)I"5�/O���t��N�2V����Q�+ϲ��)D�%��ڈ��NDh�mn�T��:����y(}�����~{i�lrK�c�;2dჰ!�t���[�b��8�3f�����d�����O��r����j����Y�]�Y�
��Ġ��l����?\�߭�d�����7�+����'ѡIU��4m��,搜: i�Z�0<Ф������x���n�x�|�?+>c��Cf������@d�8��b��	-- 3�w�&{��F
��@��O��>	�4��d�6l���`2�b���G�c�o�]{ׇ�s�b�*���2�х׳2�7L�����s�wE��h�b��T��z&�YT�//�!����sD�3��Dk���h�r�a�H9�ykP�߲PϿS~��k���́g�7ښ˟A�����1H����ˆ�
S�:m̭J*��t�����ݑ �$�]G鵭�ڝ��d�5�{W�ã��*��/wv�{�x8��" 'I��
�70
	<l�c�I>4�\duu�\G0)�gn�u�����X��j��Hn"���pcB����uݾ��v�
������)�ˊ��ކ0V���yl� JyY�$���7�2׻{#P^%�kQ=�~��N�5?"[nr�0I��Ӊ�Q��-Ȝ1��� 3����������`(�
ך��c�C0���6<ZYu��k����O�)N��k�v\�Eų�t^!���$
(��z�I�ć��:'8p�dO
�%пD։�,S^Q��K��ܠ��Y˲O�����qr�mmS2F�6Ezi�s|�40x�7��e�b	;=5(� )y�,��w>o�3�m�\8L���p�E&č:lץFУ�����nՑ����qT��3I�z6��ovd!ͬ��EJ`0CVS��z�g�F��\(��4�V^�f���������r��?g�Қo�=%R,�;]B#����O�a+���pltp�E���@c����8�F�mb(���=�;S&M����l�t�ɞ�����H��E��5#�����#x2,�rޱ~��14�_�P?}�2�3�ˈ�jm["��3v�/{3s���Y����쬗���Y76�[���uY���H��@Y�\�b��<��䲦MCᠬ����8��H!��j�6�*q��4�f�,�be�g%�(��]��E���+�e�u��˙Q�՛�;z��3Rg�Y�K(�?$�ۏ��[��[e%!r�J!! Z#Q����IA�I		I	�-B��L.j�[�;gɍ;�v����9��z��ka�Ɔ!����p�%��8P?K�/¬X�~�D��B�2�t�-�^�n�=��Sٞ�I���\3�c��+*GGR��^oW�w_ȅQ��-;7{W��t�L�%�ޒ	%{�DG���<��Y)���!�U~�z��޷D�BϠ����m��n�T�fl�	tѻn���My��y�8�hx^�U,{�Z����oAI'RP��$��]�T �@e�ӹ���c�i	��dIhA��$	)���� ����	�pŸ#�C��ٍ׌�f?wK�{���x�.-��X@��v��oM�������LV!~.v	�o�ޯ4�ws��-�ݏ��;�0/sXD��
$�O�S_�-QX�_�~G�Ðpģ$1���)Ƌ`�̍��D�gÉ���Zx��G4�Fǀ��'���Vh�%�S�"'/N���p�qU��/�u�>�U����Z_��P���
qϋ��x�!t�8�X��$ɛ(Y�wrz6��ncO�^"���B�O������J�m��X���br�g=�N�d�t�v��-.�0|�|+���(y��5���W�X $! �@���!IB[�p� ��� BB	kH�� @8B B@��H @� 0��#$�$��I!M!F!XO���U�=�����sh@�*e;2v%�JwZ�����rL��/1�f銶�H�������|�*R�gؿ9-����\P��錹no���ά�b$%�����d�L^$�ܩ:\���{|�L�#���A��eG��l@�ac9���B^�k^��tM�� U���K��ơ�X��Z\/;5�Z�����jT�Wc�C6�$`���Ssܜ�s�*d]�}�����p���j�4L��vt�^a�8�D��2-��6����$,�}X�K:	�_�-�H."q��
Dd%� l6�b������)v��jّ�R����9�r��^7���p��6�7�f�aP��K�N�`���ݼ��!-;HNC GX��~�
\Y8�G�/[�o��řyhB��%�`g�}U�]CÄ�wӸ�݀u��-�1��V\��\,�aҜ�-z[�v�ٓ�҃ŶD���J^X���WNC�L�Ffc� ���,�R�����9�W��z�������L�KY���C�V�[�� ��?��i=vف����\�dj��a�r��whR�.V����̶�p:]��.Ŕ5��Wg���SN�Pۋa]f.W\�m��USF
�,o���wBH6$$�QD#cMq��b�W	�3���o3���W`.��>�YE���4�(1��E���i!��y�3(p6��egC��T�愇��	���I5�m�#�ȊJ0���P��BX�$3�2���X��13�� |q�"Ss5�A3�~��SY���7Iˑ��=\�ͮ�{qo�ל]���d)��<G��=ג��!vfb�O�x �L��*��O�W׼]��gt���ڍt���E߼�MI �WM��H��Y3E��;3 F= ��Y��	����X<E���g�=s0`4�_P�A8��(�����U�g�>I�����X������Kt61�0 ������!�=�]|H-Ug��L�����SbߗW��<	$Y�P$��c�p��zc�3^"xmS #i��xx� �&����]��U'��4ځ"`b4�b[��gM�ConN|� �	9NI��1BZ@om��a�1w�O/wQ47ˉ��q;��Sy�'�� ��6tVbh�%�aܣ����;�08�L���_��L_}�q1c�B!�vG�OOɹ�y`K�i6ñ�&�gJ���%W�K"x�����(s���.�ݵ�eV^`�t��(X�s�`FN��H�{�G����7�QK@��D #$L�ZK�Ǖ�\S��v�&����Mfj	����Q���x�'^}�.�"��X滪�ל���ђ�A� a�v�K|F��<��mD3n�̻���×g%�3��dݛu6I�ũ���5P펓É�Wj�Ϲ*���f\ۥ�Ι�%�To҄��`��?�M�_v�qv���Ǜ"�I$�� O��{���˦���{��;�Jh��{I�<��暉�0u��@��@$$T	�Y �����:��zt�������]!00K�?U.�>xy��^��Ϝ��Ϫl�hC]�rV͗L�4y�A܈���9	z]��]��1&Z�wH����g��e��	`����mF$�x�����P�qJ:P��&�ʁ3�pV�9FvJ��c\|�M��[��A��s�ުh =���<�ܤ'�s��eCRGZ�	�(Y�d��T%�H�s�l��oq�q��C�_V�g��s��[a���%��J�j���B�g=��J5"��
h<7��膢+��O-U�g5��ր�>��p�n"��MBCE@���+��7$/n�|��{��n���]K6��0V�\�;M�����w����'.ʞ4^�i��R��[3)�3\!ufE�VU�Z�3����'9=��$�<@���[e�D#)��KɈ��F[ O&cm��?~���wi����f���%�l�B��M�8y��5x�?O�Q{���G!��mݻifH�V�j�9*����wܼ���_b]���I�]�cL�(�S�e�޽�o}�.��B�g��4�`�IO|�����V/����|eA���6�����b"B�`��p)�>���R��ř����sؠ�hۚ�z��0�������	`<+i�ټ��3��;3�Y�X#k�ۃ"��P�<�*�.�f�]/��JhR����,$����$�xt|t����� %WWh���ֱ�Z�ԁ_�q�ڶ����%��yyш�i��aƧ�n�UT$,G����r�(y��GNY
|��*�#��,x{��p�fD;[3z!���_3���C�h�'�8p�R�񹃸�JE[T�?RfL��:�t��7yzN<��{Yb�Ǹ�j^b�J�`��V��ތ����,>�F���|	s��A�"4�"H�$# �!P� �!!Q�%z����{�(04�Ѻ�ܲ.���s���B�K!ն�C��5�ͧd�>b��ۊ{��"=(b~��FS���1߽��#��A�%��I��(�$i�a�D�������MY�%㢚��M�OS�p�����l�B�<���5�$�� n����-j�b�b���↳��\f��������{����g�J�2�U-�6����(�>{f>�k�����cՊ�3S��9��MwC���܍��r�	W&�~��ܩ�=0,��߿�7O1H6�����w%��DlWL�h����a�/�6�p�ª�I,o�,7�\9ܒ�|��H���W<aL|V�3��9vr\D%W�݆ �V�YlAk��K��r/���3�g��rQk��gb��)�-� ����X:�����9!!�E����ֹ�8�}Gi�9A@�*a�:@�KJd��I$�=j(��� P�=�"��<������d�/��f�6��X�E�����c��8��k1a���b������;@�X�B �@;�X,�S �!QR�)���h#h�D �"Dh�%��튀bZ%ARD		$�I	hUgK�W� ��	 1b�EJ�؈p�X*����CXk��h�X��"QhR�f � ��6eIP�&(��*(��9���*  �A�D���40tM��`����RZ�����n��.�ل"m�)@i@iגI(>�;�׹��I ��E�0��XP�q�Н��~��5ӧ�Ӄ
����ֵ!�Gu��a�~6��wҭ�Ӛ��-�=~��8~�'�/����o#�m,!q4xtǺCC&���O?O�q�� oD�{��#��S�Ą����ӯ��w&-�l������l>����߂}��K��P'���"��_�>)��V�����H���W��*��`���aEI(�P}Jd}4�,M�v_��S9�أ����p@{�ƉW�pLƓ����K���@�0R�PN����3��d��/�����DTM�����$��u����:����H�;GcYt����
�T�ɃD�.Cq>}�ȹ9 g6^�uav�D�|Jʹ���r���+t�}q���i�dE������n)��7Y��8b-�����f����=�K�/�IG�k},o���ͽZ�'����ov�F�vZ�]�7
K'�"�D`$Tb1a���D1Q�U�"��A(��@/��S�\EA�C�Ph�Y��+ 0`�*E�� D"Db� ��F�X�DddI� $�T�DD$D@��$$�$`0E`@H� AB@� H�d)��8�@�d�	f�`�(2kXͨ�(�}@�`��ݹ�r>�'#t�j,���Q;GE l F[�jh�H�~,ǀ�n=\9�p�P�pz���AP9~��c�m��2�:������{�
8(�p4���0��$?/�i���ҵ��`"���z.�D�R�� ^�L��`�-�O��D�(F.��XX�bУ��R�BxF�o���#�#D9�o��=;��Rh<�>����`���B���k��.B�I���7���9V�tҍ�Wr�i�N uk�Lݤ�!�@p9����p�!" � � #`@9ר��V�64��>O��;jr<jY
�݃��Y̨�z�6H�"خ�抈�L���"�x���  ���좨�C[��6�1�*�_�X�4���4=>�%螯}U��[���Z��`Q���0 E�L�B���;ҕ�
��g�%$H��fA�~���<C >��c�}� �A!tB܋�*!CIT�5.�%�,���(�->A��UPЁ�+ʒ����F���cȩp>��C��/�`�$#ku��(8�("��b��v�����鬐蕅.��Ns�6�LE��v�SO#ED��g�(@�{�,W��N �� \����Rc�2f^'���C۱Ӵ���̡i�H\��X�B9���!�Z�<�R��|���n�({�=�s`��(�ǘ�o�N���n�v���|��zˢ*'�:���u5��^����Q�$�ǿ�e)�L�L�@>qED�ߌ1�eP��qt��N���'�Ǳ8��έ=g� U\ƭW!�^a��-U�;u�MؤB0���0BǠ��r���4Pr�
�p�؉`�0w�������;)�t`��2>����sT.p@�b��a^��HP�[.I��hٶ���I���,ߩ�ݓ���H��w��p�������������� Bc��Kک��BX�r��e��Sܝi+�i��8��ɧ!�p��|9Y��HȂ4�lm���+4\�.vC��C�r�W��.!���:�o&���`lD݆��`'4F(�'��J4���0{����.x�p0#�T�Yg�)�<Ơ����Q9��@T�a�d턣��c���xd�I�+�gM���;?8m���9'C�J>��C�.w��S�Z8w�@6��w$S�	r�B0